* Amplifier
.OPTIONS LIST NODE POST 
.OP 
.PRINT DC I(Rout)  I(M3)
.DC Vin 0 3 0.01

* level 1 models
.MODEL MODP PMOS LEVEL=1 VTO=-0.5 UO=500 COX=0.3e-4 LAMBDA=0.05
.MODEL MODN NMOS LEVEL=1 VTO=0.5 UO=1500 COX=0.3e-4 LAMBDA=0.05 GAMMA=0.3

VDD 9 0 DC 3
Vin 10 0 DC 1

Rin 10 11 100

Rout 16 0 1000

Vb1 12 0 DC 1

M1   13 13 9   9   MODP W=30e-6 L=0.35e-6
M2   16 12 13 13 MODP W=60e-6 L=0.35e-6
M3   16 12 14 0   MODN W=20e-6 L=0.35e-6
M4   14 11 0   0   MODN W=10e-6 L=0.35e-6

.END