* diftest
.OPTIONS LIST NODE POST 
.OP 
.PRINT DC I(M1)  I(M2)  I(D1)  I(D2)
.DC Vin 1 2 0.01
. TEMP 27

* level 1 models
.MODEL MODN1 NMOS LEVEL=1 VTO=0.5 UO=300 COX=6e-3 LAMBDA=0.05 GAMMA=0.01
.MODEL MODN2 NMOS LEVEL=1 VTO=0.3 UO=300 COX=6e-3 LAMBDA=0.05 GAMMA=0.01
.MODEL MODP1 PMOS LEVEL=1 VTO=-0.5 UO=100 COX=6e-3 LAMBDA=0.05 GAMMA=0.01
.MODEL MODP2 PMOS LEVEL=1 VTO=-0.3 UO=100 COX=6e-3 LAMBDA=0.05 GAMMA=0.01

* diode models
.MODEL DIODE D LEVEL=1 IS=1e-5

*
VDD 101 0 DC 2
Vb 111 0 DC 1
Rload1 104 0 1e5
Rload2 105 0 5

* mosfet
M1 102 112 121 0     MODN2 W=30e-6 L=0.5e-6
M2 103 112 121 0     MODN1 W=30e-6 L=0.5e-6
M3 102 111 101 101 MODP2 W=30e-6  L=0.5e-6
M4 103 111 101 101 MODP1 W=30e-6  L=0.5e-6

* diode 
D1 104 102 DIODE
D2 103 105 DIODE

* input 
VIN 112 0 1.5V
Iref 121 0 0.001

RSS 121 0 1e5


.END