*double balanced mixer
.OPTIONS LIST NODE POST 
.OP 
.ac DEC 10 0 10000000000MEG

* level 1 models
.MODEL MODP PMOS LEVEL=1 VTO=-0.58281 UO=122.4952 COX=6.058e-3 LAMBDA=0.05 CJ=4.0e-14 CAPOP=2
.MODEL MODN NMOS LEVEL=1 VTO=0.386 UO=302.38 COX=6.058e-3 LAMBDA=0.05  CJ=4.0e-14 CAPOP=2

Vdd      101 0     3V
Rload1 101 102 300
Rload2 101 103 300

* mosfets
M1 102 104 107 0 MODN W=30e-6 L=0.25e-6
M2 103 106 107 0 MODN W=30e-6 L=0.25e-6
M3 102 106 108 0 MODN W=30e-6 L=0.25e-6
M4 103 104 108 0 MODN W=30e-6 L=0.25e-6

M5 107 110 114 0 MODN W=30e-6 L=0.25e-6
M6 108 111 115 0 MODN W=30e-6 L=0.25e-6

*source degeneration
Lde1 114 129 1e-9
Rloss1 129 109 1.2
Lde2 115 139 1e-9
Rloss2 139 109 1.2

* LC tank 
Lde3 109 149 3e-9
Rloss3 149 0 3.6
Cde  109 0 9.2e-12 

*input
* SIN DC AC Freq td theta phase
Vlo+ 154 0 DC=1 AC=1,90
Rlo1 154 104 50
Vlo- 164 0 DC=1 AC=1,90
Rlo2 164 106 50

Vrf1+ 112 212 SIN 0.6 0.01 800e6 0 0 180
Vrf2+ 212 0     SIN 0    0.01 600e6 0 0 180
Vrf1- 113 213  SIN 0.6 0.01 800e6 0 0 0
Vrf2- 213 0      SIN 0    0.01 600e6 0 0 0

Rs1 112 110 25
Rs2 113 111 25

.end