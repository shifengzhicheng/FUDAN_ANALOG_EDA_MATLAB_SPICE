* RC
.OPTIONS LIST NODE POST 
.OP 
*.PRINT AC I1(M1) I2(M1) I(M2)  I(M3)  I(M4) I(Rin) I(R2) I(R3) 
.pz V(21) Vin
*.AC DEC 10 10 1e18MEG

* level 1 model
.MODEL MODN NMOS LEVEL=1 VTO=0.5 UO=1500 COX=0.3e-4 LAMBDA=0.05 Cj=4.0e-14 CAPOP=2

Vin 11 0 DC=1 AC=1,0
VDD 31 0 3
Rin 11 21 10

M1 32 21 33 0 MODN W=20e-6 L=0.35e-6

Rout 31 32 1000
Rs 33 0 10

.end
