* bjt amplifier circuit
.OPTIONS LIST NODE POST 
.OP 

Vcc 101 0 dc 9
Vbb 102 0 dc 4.0
R1 103 0 1.0e4
R2 101 104 0.2e4
R3 105 0 0.9e4
R4 101 106 1.0e4
R5 107 0 1.0e4
R6 101 108 1.0e4
Rb1 102 109 2.8e6
Rb2 108 110 1.9e5
Rb3 105 111 5.4e6

* bjt

Q1 103 109 108 MOD1
Q2 105 110 104 MOD1
Q3 107 111 106 MOD1

.MODEL MOD1 PNP IS = 2e-16 BF=100 CJE= 1e-11 CJC= 0.5e-11

.end