* RC
.OPTIONS LIST NODE POST 
.OP 
.pz V(3) Vin

Vin 1 0 AC 1

R1 1 2 10
C1 2 0 4e-6

R2 2 3 20
C2 3 0 7e-8

R3 3 4 1000
C3 3 4 5e-12

C4 4 0 8e-10

.end
