* non-inverting buffer
.OPTIONS LIST NODE POST 
.OP 
.PRINT TRAN I1(M1) I2(M1) I(M2)  I(M3)  I(M4) I(Rin) I(R2) I(R3) I(C1)
.tran 1e-9s 2e-7s

* level 1 models
.MODEL MODP PMOS LEVEL=1 VTO=-0.75 UO=500 COX=0.3e-4 LAMBDA=0.05 CJ=4.0e-14 CAPOP=0
.MODEL MODN NMOS LEVEL=1 VTO=0.83 UO=1500 COX=0.3e-4 LAMBDA=0.05 CJ=4.0e-14 CAPOP=0

VDD 103 0 3V
Vin 101 0 SIN 1.5 2 10e6 0
Rin 101 102 10

M1 107 102 103 103 MODP W=30e-6 L=0.35e-6
M2 107 102  0     0    MODN W=10e-6 L=0.35e-6
M3 104 107 103 103 MODP W=60e-6 L=0.35e-6
M4 104 107  0     0     MODN W=20e-6 L=0.35e-6

C1 104 0 0.1e-12
R2 104 115 25
L1 115 116 0.5e-12
C2 116 0 0.5e-12
R3 116 117 35
L2 117 118 0.5e-12
C3 118 0 1e-12

.END